

interface debug_intf (input clk,rst_n);

   
   


     logic debug_req_i;
     logic debug_havereset_o;
     logic debug_running_o;
     logic debug_halted_o;



endinterface : debug_intf