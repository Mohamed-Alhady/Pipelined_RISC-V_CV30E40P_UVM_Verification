class driver_config extends uvm_object ;
	
	`uvm_object_utils(driver_config)

		function  new( string name = "driver_config");
			super.new(name);
		endfunction 
endclass : driver_config

